/* Axelou Olympia
 * oaxelou@uth.gr
 * 2161
 *
 * ce430
 * Project3: VGA Controller
 *
 * Part A: VRAM Implementation
 *
 *
 * bram: Takes as input the selected address and gives as
 * output the RGB color (3bit).
 *
 * input :  clk, reset, en, address
 * output: red_output, green_output, blue_output
 *
 * Implementation:
 *   -> 3 instantiations of 16x1 Single Port BRAMs of whome we only use
 *      the 192x96 bits (12288 bits out of 16384), one for each color
 */

module bram(clk, reset, en, address, red_output, green_output, blue_output);
input clk, reset, en;
input [13:0] address;
output red_output, green_output, blue_output;

   RAMB16_S1 #(
      .INIT(1'b1),
      .SRVAL(1'b1),
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

		.INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      // the red one
      .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_2D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_2B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_2A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_29(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_27(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_26(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_24(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      // the green color
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_21(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_18(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      // the blue color
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0C(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

      // the multicolor area
      .INIT_0B(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_0A(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_09(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_08(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_07(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_06(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_05(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_04(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_03(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_02(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_01(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
      .INIT_00(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1_E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1)
    ) RED_RAMB16_S1_inst (
      .DO(red_output),
      .ADDR(address),
      .CLK(clk),
      .DI(1'b0),
      .EN(en),
      .SSR(reset),
      .WE(1'b0)
   );

   // **************************** GREEN COLOR *********************************

  RAMB16_S1 #(
    .INIT(1'b0),
    .SRVAL(1'b0),
    .WRITE_MODE("READ_FIRST"),

	  .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    // the red one
    .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2D(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_2B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_29(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_27(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_26(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_24(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    // the green color
    .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    // the blue color
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

    // the multicolor area
    .INIT_0B(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_0A(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_09(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_08(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_07(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_06(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_05(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_04(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_03(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_02(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_01(256'h99999999999999999999999999999999_99999999999999999999999999999999),
    .INIT_00(256'h99999999999999999999999999999999_99999999999999999999999999999999)
    ) GREEN_RAMB16_S1_inst (
      .DO(green_output),
      .ADDR(address),
      .CLK(clk),
      .DI(1'b0),
      .EN(en),
      .SSR(reset),
      .WE(1'b0)
      );

  // ******************************* BLUE COLOR ********************************

  RAMB16_S1 #(
     .INIT(1'b0),
     .SRVAL(1'b0),
     .WRITE_MODE("READ_FIRST"),


	  .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     // the red one
     .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_2D(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_2B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_2A(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_29(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_27(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_26(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_24(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     // the green color
     .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_21(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_1E(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_1B(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),
     .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_18(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     // the blue color
     .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
     .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),

     // the multicolor area
     .INIT_0B(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_0A(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_09(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_08(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_07(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_06(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_05(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_04(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_03(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_02(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_01(256'h87878787878787878787878787878787_87878787878787878787878787878787),
     .INIT_00(256'h87878787878787878787878787878787_87878787878787878787878787878787)
    ) BLUE_RAMB16_S1_inst (
     .DO(blue_output),
     .ADDR(address),
     .CLK(clk),
     .DI(1'b0),
     .EN(en),
     .SSR(reset),
     .WE(1'b0)
  );

endmodule
